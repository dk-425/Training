// sm_transfer_system.v

// Generated using ACDS version 22.1 922

`timescale 1 ps / 1 ps
module sm_transfer_system (
		input  wire [3:0]  buttons_export,                     //      buttons.export
		input  wire        clk_clk,                            //          clk.clk
		output wire [17:0] ext_mem_bus_tcm_address_out,        //  ext_mem_bus.tcm_address_out
		output wire [1:0]  ext_mem_bus_tcm_byteenable_n_out,   //             .tcm_byteenable_n_out
		output wire [0:0]  ext_mem_bus_tcm_outputenable_n_out, //             .tcm_outputenable_n_out
		output wire [0:0]  ext_mem_bus_tcm_write_n_out,        //             .tcm_write_n_out
		inout  wire [15:0] ext_mem_bus_tcm_data_out,           //             .tcm_data_out
		output wire [0:0]  ext_mem_bus_tcm_chipselect_n_out,   //             .tcm_chipselect_n_out
		output wire [7:0]  greenled_out_export,                // greenled_out.export
		output wire [6:0]  hex0_out_export,                    //     hex0_out.export
		output wire [6:0]  hex1_out_export,                    //     hex1_out.export
		output wire [6:0]  hex2_out_export,                    //     hex2_out.export
		output wire [6:0]  hex3_out_export,                    //     hex3_out.export
		output wire [9:0]  redled_out_export,                  //   redled_out.export
		input  wire        reset_reset_n,                      //        reset.reset_n
		output wire        ssram_clk,                          //        ssram.clk
		input  wire [9:0]  switches_export                     //     switches.export
	);

	wire         pll_outclk0_clk;                                                     // pll:outclk_0 -> [J2A_master:clk_clk, av_sm_master:clk, avalon_st_adapter:in_clk_0_clk, button_switch:csi_clock_clk, dma_source_to_ssram:clk, dma_ssram_to_led:clk, ext_mem_bus:clk, led_fifo:wrclock, led_out:csi_clock_clk, mm_interconnect_0:pll_outclk0_clk, mm_interconnect_1:pll_outclk0_clk, mm_interconnect_2:pll_outclk0_clk, reset_debounce:csi_clock_clk, rst_controller:clk, source:clk, sram_controller:clk_clk, test_mem:clk]
	wire         reset_debounce_button_qual_reset;                                    // reset_debounce:button_qual -> [J2A_master:clk_reset_reset, led_out:rsi_reset_n, mm_interconnect_0:J2A_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:led_out_reset_reset_bridge_in_reset_reset, rst_controller:reset_in0]
	wire         sram_controller_tcm_data_outen;                                      // sram_controller:tcm_data_outen -> ext_mem_bus:tcs_tcm_data_outen
	wire         sram_controller_tcm_outputenable_n_out;                              // sram_controller:tcm_outputenable_n_out -> ext_mem_bus:tcs_tcm_outputenable_n_out
	wire         sram_controller_tcm_request;                                         // sram_controller:tcm_request -> ext_mem_bus:request
	wire   [1:0] sram_controller_tcm_byteenable_n_out;                                // sram_controller:tcm_byteenable_n_out -> ext_mem_bus:tcs_tcm_byteenable_n_out
	wire         sram_controller_tcm_write_n_out;                                     // sram_controller:tcm_write_n_out -> ext_mem_bus:tcs_tcm_write_n_out
	wire         sram_controller_tcm_grant;                                           // ext_mem_bus:grant -> sram_controller:tcm_grant
	wire         sram_controller_tcm_chipselect_n_out;                                // sram_controller:tcm_chipselect_n_out -> ext_mem_bus:tcs_tcm_chipselect_n_out
	wire  [17:0] sram_controller_tcm_address_out;                                     // sram_controller:tcm_address_out -> ext_mem_bus:tcs_tcm_address_out
	wire  [15:0] sram_controller_tcm_data_out;                                        // sram_controller:tcm_data_out -> ext_mem_bus:tcs_tcm_data_out
	wire  [15:0] sram_controller_tcm_data_in;                                         // ext_mem_bus:tcs_tcm_data_in -> sram_controller:tcm_data_in
	wire         av_sm_master_avalon_master_waitrequest;                              // mm_interconnect_0:av_sm_master_avalon_master_waitrequest -> av_sm_master:am_waitreq
	wire  [31:0] av_sm_master_avalon_master_readdata;                                 // mm_interconnect_0:av_sm_master_avalon_master_readdata -> av_sm_master:am_data_in
	wire  [31:0] av_sm_master_avalon_master_address;                                  // av_sm_master:am_addr -> mm_interconnect_0:av_sm_master_avalon_master_address
	wire         av_sm_master_avalon_master_read;                                     // av_sm_master:am_rd -> mm_interconnect_0:av_sm_master_avalon_master_read
	wire  [31:0] av_sm_master_avalon_master_writedata;                                // av_sm_master:am_data_out -> mm_interconnect_0:av_sm_master_avalon_master_writedata
	wire         av_sm_master_avalon_master_write;                                    // av_sm_master:am_wr -> mm_interconnect_0:av_sm_master_avalon_master_write
	wire  [31:0] j2a_master_master_readdata;                                          // mm_interconnect_0:J2A_master_master_readdata -> J2A_master:master_readdata
	wire         j2a_master_master_waitrequest;                                       // mm_interconnect_0:J2A_master_master_waitrequest -> J2A_master:master_waitrequest
	wire  [31:0] j2a_master_master_address;                                           // J2A_master:master_address -> mm_interconnect_0:J2A_master_master_address
	wire         j2a_master_master_read;                                              // J2A_master:master_read -> mm_interconnect_0:J2A_master_master_read
	wire   [3:0] j2a_master_master_byteenable;                                        // J2A_master:master_byteenable -> mm_interconnect_0:J2A_master_master_byteenable
	wire         j2a_master_master_readdatavalid;                                     // mm_interconnect_0:J2A_master_master_readdatavalid -> J2A_master:master_readdatavalid
	wire         j2a_master_master_write;                                             // J2A_master:master_write -> mm_interconnect_0:J2A_master_master_write
	wire  [31:0] j2a_master_master_writedata;                                         // J2A_master:master_writedata -> mm_interconnect_0:J2A_master_master_writedata
	wire  [31:0] led_out_swpb_readdata;                                               // mm_interconnect_0:led_out_swpb_readdata -> led_out:avm_swpb_readdata
	wire         led_out_swpb_waitrequest;                                            // mm_interconnect_0:led_out_swpb_waitrequest -> led_out:avm_swpb_waitrequest
	wire  [31:0] led_out_swpb_address;                                                // led_out:avm_swpb_address -> mm_interconnect_0:led_out_swpb_address
	wire         led_out_swpb_read;                                                   // led_out:avm_swpb_read_n -> mm_interconnect_0:led_out_swpb_read
	wire         dma_ssram_to_led_write_master_chipselect;                            // dma_ssram_to_led:write_chipselect -> mm_interconnect_0:dma_ssram_to_led_write_master_chipselect
	wire         dma_ssram_to_led_write_master_waitrequest;                           // mm_interconnect_0:dma_ssram_to_led_write_master_waitrequest -> dma_ssram_to_led:write_waitrequest
	wire  [20:0] dma_ssram_to_led_write_master_address;                               // dma_ssram_to_led:write_address -> mm_interconnect_0:dma_ssram_to_led_write_master_address
	wire   [3:0] dma_ssram_to_led_write_master_byteenable;                            // dma_ssram_to_led:write_byteenable -> mm_interconnect_0:dma_ssram_to_led_write_master_byteenable
	wire         dma_ssram_to_led_write_master_write;                                 // dma_ssram_to_led:write_write_n -> mm_interconnect_0:dma_ssram_to_led_write_master_write
	wire  [31:0] dma_ssram_to_led_write_master_writedata;                             // dma_ssram_to_led:write_writedata -> mm_interconnect_0:dma_ssram_to_led_write_master_writedata
	wire  [31:0] mm_interconnect_0_button_switch_buttonreg_readdata;                  // button_switch:avs_buttonreg_readdata -> mm_interconnect_0:button_switch_buttonreg_readdata
	wire   [1:0] mm_interconnect_0_button_switch_buttonreg_address;                   // mm_interconnect_0:button_switch_buttonreg_address -> button_switch:avs_buttonreg_address
	wire         mm_interconnect_0_button_switch_buttonreg_read;                      // mm_interconnect_0:button_switch_buttonreg_read -> button_switch:avs_buttonreg_read
	wire         mm_interconnect_0_button_switch_buttonreg_write;                     // mm_interconnect_0:button_switch_buttonreg_write -> button_switch:avs_buttonreg_write
	wire  [31:0] mm_interconnect_0_button_switch_buttonreg_writedata;                 // mm_interconnect_0:button_switch_buttonreg_writedata -> button_switch:avs_buttonreg_writedata
	wire         mm_interconnect_0_dma_ssram_to_led_control_port_slave_chipselect;    // mm_interconnect_0:dma_ssram_to_led_control_port_slave_chipselect -> dma_ssram_to_led:dma_ctl_chipselect
	wire  [20:0] mm_interconnect_0_dma_ssram_to_led_control_port_slave_readdata;      // dma_ssram_to_led:dma_ctl_readdata -> mm_interconnect_0:dma_ssram_to_led_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_dma_ssram_to_led_control_port_slave_address;       // mm_interconnect_0:dma_ssram_to_led_control_port_slave_address -> dma_ssram_to_led:dma_ctl_address
	wire         mm_interconnect_0_dma_ssram_to_led_control_port_slave_write;         // mm_interconnect_0:dma_ssram_to_led_control_port_slave_write -> dma_ssram_to_led:dma_ctl_write_n
	wire  [20:0] mm_interconnect_0_dma_ssram_to_led_control_port_slave_writedata;     // mm_interconnect_0:dma_ssram_to_led_control_port_slave_writedata -> dma_ssram_to_led:dma_ctl_writedata
	wire         mm_interconnect_0_dma_source_to_ssram_control_port_slave_chipselect; // mm_interconnect_0:dma_source_to_ssram_control_port_slave_chipselect -> dma_source_to_ssram:dma_ctl_chipselect
	wire  [17:0] mm_interconnect_0_dma_source_to_ssram_control_port_slave_readdata;   // dma_source_to_ssram:dma_ctl_readdata -> mm_interconnect_0:dma_source_to_ssram_control_port_slave_readdata
	wire   [2:0] mm_interconnect_0_dma_source_to_ssram_control_port_slave_address;    // mm_interconnect_0:dma_source_to_ssram_control_port_slave_address -> dma_source_to_ssram:dma_ctl_address
	wire         mm_interconnect_0_dma_source_to_ssram_control_port_slave_write;      // mm_interconnect_0:dma_source_to_ssram_control_port_slave_write -> dma_source_to_ssram:dma_ctl_write_n
	wire  [17:0] mm_interconnect_0_dma_source_to_ssram_control_port_slave_writedata;  // mm_interconnect_0:dma_source_to_ssram_control_port_slave_writedata -> dma_source_to_ssram:dma_ctl_writedata
	wire         mm_interconnect_0_led_fifo_in_waitrequest;                           // led_fifo:avalonmm_write_slave_waitrequest -> mm_interconnect_0:led_fifo_in_waitrequest
	wire   [0:0] mm_interconnect_0_led_fifo_in_address;                               // mm_interconnect_0:led_fifo_in_address -> led_fifo:avalonmm_write_slave_address
	wire         mm_interconnect_0_led_fifo_in_write;                                 // mm_interconnect_0:led_fifo_in_write -> led_fifo:avalonmm_write_slave_write
	wire  [31:0] mm_interconnect_0_led_fifo_in_writedata;                             // mm_interconnect_0:led_fifo_in_writedata -> led_fifo:avalonmm_write_slave_writedata
	wire  [31:0] mm_interconnect_0_led_out_led_readdata;                              // led_out:avs_led_readdata -> mm_interconnect_0:led_out_led_readdata
	wire   [1:0] mm_interconnect_0_led_out_led_address;                               // mm_interconnect_0:led_out_led_address -> led_out:avs_led_address
	wire         mm_interconnect_0_led_out_led_read;                                  // mm_interconnect_0:led_out_led_read -> led_out:avs_led_read
	wire         mm_interconnect_0_led_out_led_write;                                 // mm_interconnect_0:led_out_led_write -> led_out:avs_led_write
	wire  [31:0] mm_interconnect_0_led_out_led_writedata;                             // mm_interconnect_0:led_out_led_writedata -> led_out:avs_led_writedata
	wire         mm_interconnect_0_test_mem_s1_chipselect;                            // mm_interconnect_0:test_mem_s1_chipselect -> test_mem:chipselect
	wire  [31:0] mm_interconnect_0_test_mem_s1_readdata;                              // test_mem:readdata -> mm_interconnect_0:test_mem_s1_readdata
	wire  [10:0] mm_interconnect_0_test_mem_s1_address;                               // mm_interconnect_0:test_mem_s1_address -> test_mem:address
	wire   [3:0] mm_interconnect_0_test_mem_s1_byteenable;                            // mm_interconnect_0:test_mem_s1_byteenable -> test_mem:byteenable
	wire         mm_interconnect_0_test_mem_s1_write;                                 // mm_interconnect_0:test_mem_s1_write -> test_mem:write
	wire  [31:0] mm_interconnect_0_test_mem_s1_writedata;                             // mm_interconnect_0:test_mem_s1_writedata -> test_mem:writedata
	wire         mm_interconnect_0_test_mem_s1_clken;                                 // mm_interconnect_0:test_mem_s1_clken -> test_mem:clken
	wire         dma_source_to_ssram_read_master_chipselect;                          // dma_source_to_ssram:read_chipselect -> mm_interconnect_1:dma_source_to_ssram_read_master_chipselect
	wire  [31:0] dma_source_to_ssram_read_master_readdata;                            // mm_interconnect_1:dma_source_to_ssram_read_master_readdata -> dma_source_to_ssram:read_readdata
	wire         dma_source_to_ssram_read_master_waitrequest;                         // mm_interconnect_1:dma_source_to_ssram_read_master_waitrequest -> dma_source_to_ssram:read_waitrequest
	wire  [12:0] dma_source_to_ssram_read_master_address;                             // dma_source_to_ssram:read_address -> mm_interconnect_1:dma_source_to_ssram_read_master_address
	wire         dma_source_to_ssram_read_master_read;                                // dma_source_to_ssram:read_read_n -> mm_interconnect_1:dma_source_to_ssram_read_master_read
	wire         dma_source_to_ssram_read_master_readdatavalid;                       // mm_interconnect_1:dma_source_to_ssram_read_master_readdatavalid -> dma_source_to_ssram:read_readdatavalid
	wire         mm_interconnect_1_source_s1_chipselect;                              // mm_interconnect_1:source_s1_chipselect -> source:chipselect
	wire  [31:0] mm_interconnect_1_source_s1_readdata;                                // source:readdata -> mm_interconnect_1:source_s1_readdata
	wire         mm_interconnect_1_source_s1_debugaccess;                             // mm_interconnect_1:source_s1_debugaccess -> source:debugaccess
	wire  [10:0] mm_interconnect_1_source_s1_address;                                 // mm_interconnect_1:source_s1_address -> source:address
	wire   [3:0] mm_interconnect_1_source_s1_byteenable;                              // mm_interconnect_1:source_s1_byteenable -> source:byteenable
	wire         mm_interconnect_1_source_s1_write;                                   // mm_interconnect_1:source_s1_write -> source:write
	wire  [31:0] mm_interconnect_1_source_s1_writedata;                               // mm_interconnect_1:source_s1_writedata -> source:writedata
	wire         mm_interconnect_1_source_s1_clken;                                   // mm_interconnect_1:source_s1_clken -> source:clken
	wire         dma_ssram_to_led_read_master_chipselect;                             // dma_ssram_to_led:read_chipselect -> mm_interconnect_2:dma_ssram_to_led_read_master_chipselect
	wire  [31:0] dma_ssram_to_led_read_master_readdata;                               // mm_interconnect_2:dma_ssram_to_led_read_master_readdata -> dma_ssram_to_led:read_readdata
	wire         dma_ssram_to_led_read_master_waitrequest;                            // mm_interconnect_2:dma_ssram_to_led_read_master_waitrequest -> dma_ssram_to_led:read_waitrequest
	wire  [17:0] dma_ssram_to_led_read_master_address;                                // dma_ssram_to_led:read_address -> mm_interconnect_2:dma_ssram_to_led_read_master_address
	wire         dma_ssram_to_led_read_master_read;                                   // dma_ssram_to_led:read_read_n -> mm_interconnect_2:dma_ssram_to_led_read_master_read
	wire         dma_ssram_to_led_read_master_readdatavalid;                          // mm_interconnect_2:dma_ssram_to_led_read_master_readdatavalid -> dma_ssram_to_led:read_readdatavalid
	wire         dma_source_to_ssram_write_master_chipselect;                         // dma_source_to_ssram:write_chipselect -> mm_interconnect_2:dma_source_to_ssram_write_master_chipselect
	wire         dma_source_to_ssram_write_master_waitrequest;                        // mm_interconnect_2:dma_source_to_ssram_write_master_waitrequest -> dma_source_to_ssram:write_waitrequest
	wire  [17:0] dma_source_to_ssram_write_master_address;                            // dma_source_to_ssram:write_address -> mm_interconnect_2:dma_source_to_ssram_write_master_address
	wire   [3:0] dma_source_to_ssram_write_master_byteenable;                         // dma_source_to_ssram:write_byteenable -> mm_interconnect_2:dma_source_to_ssram_write_master_byteenable
	wire         dma_source_to_ssram_write_master_write;                              // dma_source_to_ssram:write_write_n -> mm_interconnect_2:dma_source_to_ssram_write_master_write
	wire  [31:0] dma_source_to_ssram_write_master_writedata;                          // dma_source_to_ssram:write_writedata -> mm_interconnect_2:dma_source_to_ssram_write_master_writedata
	wire  [15:0] mm_interconnect_2_sram_controller_uas_readdata;                      // sram_controller:uas_readdata -> mm_interconnect_2:sram_controller_uas_readdata
	wire         mm_interconnect_2_sram_controller_uas_waitrequest;                   // sram_controller:uas_waitrequest -> mm_interconnect_2:sram_controller_uas_waitrequest
	wire         mm_interconnect_2_sram_controller_uas_debugaccess;                   // mm_interconnect_2:sram_controller_uas_debugaccess -> sram_controller:uas_debugaccess
	wire  [17:0] mm_interconnect_2_sram_controller_uas_address;                       // mm_interconnect_2:sram_controller_uas_address -> sram_controller:uas_address
	wire         mm_interconnect_2_sram_controller_uas_read;                          // mm_interconnect_2:sram_controller_uas_read -> sram_controller:uas_read
	wire   [1:0] mm_interconnect_2_sram_controller_uas_byteenable;                    // mm_interconnect_2:sram_controller_uas_byteenable -> sram_controller:uas_byteenable
	wire         mm_interconnect_2_sram_controller_uas_readdatavalid;                 // sram_controller:uas_readdatavalid -> mm_interconnect_2:sram_controller_uas_readdatavalid
	wire         mm_interconnect_2_sram_controller_uas_lock;                          // mm_interconnect_2:sram_controller_uas_lock -> sram_controller:uas_lock
	wire         mm_interconnect_2_sram_controller_uas_write;                         // mm_interconnect_2:sram_controller_uas_write -> sram_controller:uas_write
	wire  [15:0] mm_interconnect_2_sram_controller_uas_writedata;                     // mm_interconnect_2:sram_controller_uas_writedata -> sram_controller:uas_writedata
	wire   [1:0] mm_interconnect_2_sram_controller_uas_burstcount;                    // mm_interconnect_2:sram_controller_uas_burstcount -> sram_controller:uas_burstcount
	wire         led_fifo_out_valid;                                                  // led_fifo:avalonst_source_valid -> avalon_st_adapter:in_0_valid
	wire  [31:0] led_fifo_out_data;                                                   // led_fifo:avalonst_source_data -> avalon_st_adapter:in_0_data
	wire         led_fifo_out_ready;                                                  // avalon_st_adapter:in_0_ready -> led_fifo:avalonst_source_ready
	wire         avalon_st_adapter_out_0_valid;                                       // avalon_st_adapter:out_0_valid -> led_out:asi_ledfifo_valid
	wire  [31:0] avalon_st_adapter_out_0_data;                                        // avalon_st_adapter:out_0_data -> led_out:asi_ledfifo_data
	wire         avalon_st_adapter_out_0_ready;                                       // led_out:asi_ledfifo_ready -> avalon_st_adapter:out_0_ready
	wire         rst_controller_reset_out_reset;                                      // rst_controller:reset_out -> [av_sm_master:rst, avalon_st_adapter:in_rst_0_reset, button_switch:rsi_reset_n, dma_source_to_ssram:system_reset_n, dma_ssram_to_led:system_reset_n, ext_mem_bus:reset, led_fifo:reset_n, mm_interconnect_0:av_sm_master_reset_reset_bridge_in_reset_reset, mm_interconnect_1:dma_source_to_ssram_reset_reset_bridge_in_reset_reset, mm_interconnect_2:dma_ssram_to_led_reset_reset_bridge_in_reset_reset, source:reset, sram_controller:reset_reset, test_mem:reset]
	wire         j2a_master_master_reset_reset;                                       // J2A_master:master_reset_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                  // rst_controller_001:reset_out -> pll:rst

	sm_transfer_system_J2A_master #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) j2a_master (
		.clk_clk              (pll_outclk0_clk),                  //          clk.clk
		.clk_reset_reset      (reset_debounce_button_qual_reset), //    clk_reset.reset
		.master_address       (j2a_master_master_address),        //       master.address
		.master_readdata      (j2a_master_master_readdata),       //             .readdata
		.master_read          (j2a_master_master_read),           //             .read
		.master_write         (j2a_master_master_write),          //             .write
		.master_writedata     (j2a_master_master_writedata),      //             .writedata
		.master_waitrequest   (j2a_master_master_waitrequest),    //             .waitrequest
		.master_readdatavalid (j2a_master_master_readdatavalid),  //             .readdatavalid
		.master_byteenable    (j2a_master_master_byteenable),     //             .byteenable
		.master_reset_reset   (j2a_master_master_reset_reset)     // master_reset.reset
	);

	avalon_state_machine_master av_sm_master (
		.clk         (pll_outclk0_clk),                        //         clock.clk
		.rst         (rst_controller_reset_out_reset),         //         reset.reset
		.am_waitreq  (av_sm_master_avalon_master_waitrequest), // avalon_master.waitrequest
		.am_data_in  (av_sm_master_avalon_master_readdata),    //              .readdata
		.am_addr     (av_sm_master_avalon_master_address),     //              .address
		.am_data_out (av_sm_master_avalon_master_writedata),   //              .writedata
		.am_rd       (av_sm_master_avalon_master_read),        //              .read
		.am_wr       (av_sm_master_avalon_master_write)        //              .write
	);

	button_switch_pio #(
		.BUTTON_WIDTH (4),
		.SWITCH_WIDTH (10)
	) button_switch (
		.csi_clock_clk           (pll_outclk0_clk),                                     //          clock.clk
		.rsi_reset_n             (~rst_controller_reset_out_reset),                     //          reset.reset_n
		.avs_buttonreg_address   (mm_interconnect_0_button_switch_buttonreg_address),   //      buttonreg.address
		.avs_buttonreg_writedata (mm_interconnect_0_button_switch_buttonreg_writedata), //               .writedata
		.avs_buttonreg_readdata  (mm_interconnect_0_button_switch_buttonreg_readdata),  //               .readdata
		.avs_buttonreg_write     (mm_interconnect_0_button_switch_buttonreg_write),     //               .write
		.avs_buttonreg_read      (mm_interconnect_0_button_switch_buttonreg_read),      //               .read
		.coe_buttons_in          (buttons_export),                                      // button_conduit.export
		.coe_switches_in         (switches_export)                                      // switch_conduit.export
	);

	sm_transfer_system_dma_source_to_ssram dma_source_to_ssram (
		.clk                (pll_outclk0_clk),                                                     //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                                     //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_dma_source_to_ssram_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_dma_source_to_ssram_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_dma_source_to_ssram_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_dma_source_to_ssram_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_dma_source_to_ssram_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (),                                                                    //                irq.irq
		.read_address       (dma_source_to_ssram_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_source_to_ssram_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_source_to_ssram_read_master_read),                                //                   .read_n
		.read_readdata      (dma_source_to_ssram_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_source_to_ssram_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_source_to_ssram_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_source_to_ssram_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_source_to_ssram_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_source_to_ssram_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_source_to_ssram_write_master_write),                              //                   .write_n
		.write_writedata    (dma_source_to_ssram_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_source_to_ssram_write_master_byteenable)                          //                   .byteenable
	);

	sm_transfer_system_dma_ssram_to_led dma_ssram_to_led (
		.clk                (pll_outclk0_clk),                                                  //                clk.clk
		.system_reset_n     (~rst_controller_reset_out_reset),                                  //              reset.reset_n
		.dma_ctl_address    (mm_interconnect_0_dma_ssram_to_led_control_port_slave_address),    // control_port_slave.address
		.dma_ctl_chipselect (mm_interconnect_0_dma_ssram_to_led_control_port_slave_chipselect), //                   .chipselect
		.dma_ctl_readdata   (mm_interconnect_0_dma_ssram_to_led_control_port_slave_readdata),   //                   .readdata
		.dma_ctl_write_n    (~mm_interconnect_0_dma_ssram_to_led_control_port_slave_write),     //                   .write_n
		.dma_ctl_writedata  (mm_interconnect_0_dma_ssram_to_led_control_port_slave_writedata),  //                   .writedata
		.dma_ctl_irq        (),                                                                 //                irq.irq
		.read_address       (dma_ssram_to_led_read_master_address),                             //        read_master.address
		.read_chipselect    (dma_ssram_to_led_read_master_chipselect),                          //                   .chipselect
		.read_read_n        (dma_ssram_to_led_read_master_read),                                //                   .read_n
		.read_readdata      (dma_ssram_to_led_read_master_readdata),                            //                   .readdata
		.read_readdatavalid (dma_ssram_to_led_read_master_readdatavalid),                       //                   .readdatavalid
		.read_waitrequest   (dma_ssram_to_led_read_master_waitrequest),                         //                   .waitrequest
		.write_address      (dma_ssram_to_led_write_master_address),                            //       write_master.address
		.write_chipselect   (dma_ssram_to_led_write_master_chipselect),                         //                   .chipselect
		.write_waitrequest  (dma_ssram_to_led_write_master_waitrequest),                        //                   .waitrequest
		.write_write_n      (dma_ssram_to_led_write_master_write),                              //                   .write_n
		.write_writedata    (dma_ssram_to_led_write_master_writedata),                          //                   .writedata
		.write_byteenable   (dma_ssram_to_led_write_master_byteenable)                          //                   .byteenable
	);

	sm_transfer_system_ext_mem_bus ext_mem_bus (
		.clk                        (pll_outclk0_clk),                        //   clk.clk
		.reset                      (rst_controller_reset_out_reset),         // reset.reset
		.request                    (sram_controller_tcm_request),            //   tcs.request
		.grant                      (sram_controller_tcm_grant),              //      .grant
		.tcs_tcm_address_out        (sram_controller_tcm_address_out),        //      .address_out
		.tcs_tcm_byteenable_n_out   (sram_controller_tcm_byteenable_n_out),   //      .byteenable_n_out
		.tcs_tcm_outputenable_n_out (sram_controller_tcm_outputenable_n_out), //      .outputenable_n_out
		.tcs_tcm_write_n_out        (sram_controller_tcm_write_n_out),        //      .write_n_out
		.tcs_tcm_data_out           (sram_controller_tcm_data_out),           //      .data_out
		.tcs_tcm_data_outen         (sram_controller_tcm_data_outen),         //      .data_outen
		.tcs_tcm_data_in            (sram_controller_tcm_data_in),            //      .data_in
		.tcs_tcm_chipselect_n_out   (sram_controller_tcm_chipselect_n_out),   //      .chipselect_n_out
		.tcm_address_out            (ext_mem_bus_tcm_address_out),            //   out.tcm_address_out
		.tcm_byteenable_n_out       (ext_mem_bus_tcm_byteenable_n_out),       //      .tcm_byteenable_n_out
		.tcm_outputenable_n_out     (ext_mem_bus_tcm_outputenable_n_out),     //      .tcm_outputenable_n_out
		.tcm_write_n_out            (ext_mem_bus_tcm_write_n_out),            //      .tcm_write_n_out
		.tcm_data_out               (ext_mem_bus_tcm_data_out),               //      .tcm_data_out
		.tcm_chipselect_n_out       (ext_mem_bus_tcm_chipselect_n_out)        //      .tcm_chipselect_n_out
	);

	sm_transfer_system_led_fifo led_fifo (
		.wrclock                          (pll_outclk0_clk),                           //   clk_in.clk
		.reset_n                          (~rst_controller_reset_out_reset),           // reset_in.reset_n
		.avalonmm_write_slave_writedata   (mm_interconnect_0_led_fifo_in_writedata),   //       in.writedata
		.avalonmm_write_slave_write       (mm_interconnect_0_led_fifo_in_write),       //         .write
		.avalonmm_write_slave_address     (mm_interconnect_0_led_fifo_in_address),     //         .address
		.avalonmm_write_slave_waitrequest (mm_interconnect_0_led_fifo_in_waitrequest), //         .waitrequest
		.avalonst_source_valid            (led_fifo_out_valid),                        //      out.valid
		.avalonst_source_data             (led_fifo_out_data),                         //         .data
		.avalonst_source_ready            (led_fifo_out_ready)                         //         .ready
	);

	avalon_st_mm_led #(
		.COUNT_MAX   (34'b0000000100111111111111111111111111),
		.GREEN_WIDTH (8),
		.RED_WIDTH   (10)
	) led_out (
		.csi_clock_clk        (pll_outclk0_clk),                         //        clock.clk
		.rsi_reset_n          (~reset_debounce_button_qual_reset),       //        reset.reset_n
		.avs_led_writedata    (mm_interconnect_0_led_out_led_writedata), //          led.writedata
		.avs_led_address      (mm_interconnect_0_led_out_led_address),   //             .address
		.avs_led_readdata     (mm_interconnect_0_led_out_led_readdata),  //             .readdata
		.avs_led_write        (mm_interconnect_0_led_out_led_write),     //             .write
		.avs_led_read         (mm_interconnect_0_led_out_led_read),      //             .read
		.avm_swpb_address     (led_out_swpb_address),                    //         swpb.address
		.avm_swpb_readdata    (led_out_swpb_readdata),                   //             .readdata
		.avm_swpb_waitrequest (led_out_swpb_waitrequest),                //             .waitrequest
		.avm_swpb_read_n      (led_out_swpb_read),                       //             .read_n
		.asi_ledfifo_valid    (avalon_st_adapter_out_0_valid),           //      ledfifo.valid
		.asi_ledfifo_data     (avalon_st_adapter_out_0_data),            //             .data
		.asi_ledfifo_ready    (avalon_st_adapter_out_0_ready),           //             .ready
		.coe_greenled_out     (greenled_out_export),                     // greenled_out.export
		.coe_hex0_out         (hex0_out_export),                         //     hex0_out.export
		.coe_redled_out       (redled_out_export),                       //   redled_out.export
		.coe_hex1_out         (hex1_out_export),                         //     hex1_out.export
		.coe_hex2_out         (hex2_out_export),                         //     hex2_out.export
		.coe_hex3_out         (hex3_out_export)                          //     hex3_out.export
	);

	sm_transfer_system_pll pll (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_001_reset_out_reset), //   reset.reset
		.outclk_0 (pll_outclk0_clk),                    // outclk0.clk
		.outclk_1 (ssram_clk),                          // outclk1.clk
		.locked   ()                                    //  locked.export
	);

	button_debounce reset_debounce (
		.csi_clock_clk (pll_outclk0_clk),                  //              clock.clk
		.coe_button_in (reset_reset_n),                    // button_debounce_in.reset_n
		.button_qual   (reset_debounce_button_qual_reset), //        button_qual.reset
		.button_qual_n ()                                  //      button_qual_n.reset_n
	);

	sm_transfer_system_source source (
		.clk         (pll_outclk0_clk),                         //   clk1.clk
		.address     (mm_interconnect_1_source_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_1_source_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_1_source_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_1_source_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_1_source_s1_write),       //       .write
		.readdata    (mm_interconnect_1_source_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_1_source_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_1_source_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),          // reset1.reset
		.reset_req   (1'b0),                                    // (terminated)
		.freeze      (1'b0)                                     // (terminated)
	);

	sm_transfer_system_sram_controller #(
		.TCM_ADDRESS_W                  (18),
		.TCM_DATA_W                     (16),
		.TCM_BYTEENABLE_W               (2),
		.TCM_READ_WAIT                  (10),
		.TCM_WRITE_WAIT                 (10),
		.TCM_SETUP_WAIT                 (10),
		.TCM_DATA_HOLD                  (10),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (2),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (0),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (1),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (1),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (0),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (1),
		.ACTIVE_LOW_OUTPUTENABLE        (1),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) sram_controller (
		.clk_clk                (pll_outclk0_clk),                                     //   clk.clk
		.reset_reset            (rst_controller_reset_out_reset),                      // reset.reset
		.uas_address            (mm_interconnect_2_sram_controller_uas_address),       //   uas.address
		.uas_burstcount         (mm_interconnect_2_sram_controller_uas_burstcount),    //      .burstcount
		.uas_read               (mm_interconnect_2_sram_controller_uas_read),          //      .read
		.uas_write              (mm_interconnect_2_sram_controller_uas_write),         //      .write
		.uas_waitrequest        (mm_interconnect_2_sram_controller_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid      (mm_interconnect_2_sram_controller_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable         (mm_interconnect_2_sram_controller_uas_byteenable),    //      .byteenable
		.uas_readdata           (mm_interconnect_2_sram_controller_uas_readdata),      //      .readdata
		.uas_writedata          (mm_interconnect_2_sram_controller_uas_writedata),     //      .writedata
		.uas_lock               (mm_interconnect_2_sram_controller_uas_lock),          //      .lock
		.uas_debugaccess        (mm_interconnect_2_sram_controller_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out        (sram_controller_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_chipselect_n_out   (sram_controller_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_outputenable_n_out (sram_controller_tcm_outputenable_n_out),              //      .outputenable_n_out
		.tcm_request            (sram_controller_tcm_request),                         //      .request
		.tcm_grant              (sram_controller_tcm_grant),                           //      .grant
		.tcm_address_out        (sram_controller_tcm_address_out),                     //      .address_out
		.tcm_byteenable_n_out   (sram_controller_tcm_byteenable_n_out),                //      .byteenable_n_out
		.tcm_data_out           (sram_controller_tcm_data_out),                        //      .data_out
		.tcm_data_outen         (sram_controller_tcm_data_outen),                      //      .data_outen
		.tcm_data_in            (sram_controller_tcm_data_in)                          //      .data_in
	);

	sm_transfer_system_test_mem test_mem (
		.clk        (pll_outclk0_clk),                          //   clk1.clk
		.address    (mm_interconnect_0_test_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_test_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_test_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_test_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_test_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_test_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_test_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),           // reset1.reset
		.reset_req  (1'b0),                                     // (terminated)
		.freeze     (1'b0)                                      // (terminated)
	);

	sm_transfer_system_mm_interconnect_0 mm_interconnect_0 (
		.pll_outclk0_clk                                   (pll_outclk0_clk),                                                     //                                pll_outclk0.clk
		.av_sm_master_reset_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                                      //   av_sm_master_reset_reset_bridge_in_reset.reset
		.J2A_master_clk_reset_reset_bridge_in_reset_reset  (reset_debounce_button_qual_reset),                                    // J2A_master_clk_reset_reset_bridge_in_reset.reset
		.led_out_reset_reset_bridge_in_reset_reset         (reset_debounce_button_qual_reset),                                    //        led_out_reset_reset_bridge_in_reset.reset
		.av_sm_master_avalon_master_address                (av_sm_master_avalon_master_address),                                  //                 av_sm_master_avalon_master.address
		.av_sm_master_avalon_master_waitrequest            (av_sm_master_avalon_master_waitrequest),                              //                                           .waitrequest
		.av_sm_master_avalon_master_read                   (av_sm_master_avalon_master_read),                                     //                                           .read
		.av_sm_master_avalon_master_readdata               (av_sm_master_avalon_master_readdata),                                 //                                           .readdata
		.av_sm_master_avalon_master_write                  (av_sm_master_avalon_master_write),                                    //                                           .write
		.av_sm_master_avalon_master_writedata              (av_sm_master_avalon_master_writedata),                                //                                           .writedata
		.dma_ssram_to_led_write_master_address             (dma_ssram_to_led_write_master_address),                               //              dma_ssram_to_led_write_master.address
		.dma_ssram_to_led_write_master_waitrequest         (dma_ssram_to_led_write_master_waitrequest),                           //                                           .waitrequest
		.dma_ssram_to_led_write_master_byteenable          (dma_ssram_to_led_write_master_byteenable),                            //                                           .byteenable
		.dma_ssram_to_led_write_master_chipselect          (dma_ssram_to_led_write_master_chipselect),                            //                                           .chipselect
		.dma_ssram_to_led_write_master_write               (~dma_ssram_to_led_write_master_write),                                //                                           .write
		.dma_ssram_to_led_write_master_writedata           (dma_ssram_to_led_write_master_writedata),                             //                                           .writedata
		.J2A_master_master_address                         (j2a_master_master_address),                                           //                          J2A_master_master.address
		.J2A_master_master_waitrequest                     (j2a_master_master_waitrequest),                                       //                                           .waitrequest
		.J2A_master_master_byteenable                      (j2a_master_master_byteenable),                                        //                                           .byteenable
		.J2A_master_master_read                            (j2a_master_master_read),                                              //                                           .read
		.J2A_master_master_readdata                        (j2a_master_master_readdata),                                          //                                           .readdata
		.J2A_master_master_readdatavalid                   (j2a_master_master_readdatavalid),                                     //                                           .readdatavalid
		.J2A_master_master_write                           (j2a_master_master_write),                                             //                                           .write
		.J2A_master_master_writedata                       (j2a_master_master_writedata),                                         //                                           .writedata
		.led_out_swpb_address                              (led_out_swpb_address),                                                //                               led_out_swpb.address
		.led_out_swpb_waitrequest                          (led_out_swpb_waitrequest),                                            //                                           .waitrequest
		.led_out_swpb_read                                 (~led_out_swpb_read),                                                  //                                           .read
		.led_out_swpb_readdata                             (led_out_swpb_readdata),                                               //                                           .readdata
		.button_switch_buttonreg_address                   (mm_interconnect_0_button_switch_buttonreg_address),                   //                    button_switch_buttonreg.address
		.button_switch_buttonreg_write                     (mm_interconnect_0_button_switch_buttonreg_write),                     //                                           .write
		.button_switch_buttonreg_read                      (mm_interconnect_0_button_switch_buttonreg_read),                      //                                           .read
		.button_switch_buttonreg_readdata                  (mm_interconnect_0_button_switch_buttonreg_readdata),                  //                                           .readdata
		.button_switch_buttonreg_writedata                 (mm_interconnect_0_button_switch_buttonreg_writedata),                 //                                           .writedata
		.dma_source_to_ssram_control_port_slave_address    (mm_interconnect_0_dma_source_to_ssram_control_port_slave_address),    //     dma_source_to_ssram_control_port_slave.address
		.dma_source_to_ssram_control_port_slave_write      (mm_interconnect_0_dma_source_to_ssram_control_port_slave_write),      //                                           .write
		.dma_source_to_ssram_control_port_slave_readdata   (mm_interconnect_0_dma_source_to_ssram_control_port_slave_readdata),   //                                           .readdata
		.dma_source_to_ssram_control_port_slave_writedata  (mm_interconnect_0_dma_source_to_ssram_control_port_slave_writedata),  //                                           .writedata
		.dma_source_to_ssram_control_port_slave_chipselect (mm_interconnect_0_dma_source_to_ssram_control_port_slave_chipselect), //                                           .chipselect
		.dma_ssram_to_led_control_port_slave_address       (mm_interconnect_0_dma_ssram_to_led_control_port_slave_address),       //        dma_ssram_to_led_control_port_slave.address
		.dma_ssram_to_led_control_port_slave_write         (mm_interconnect_0_dma_ssram_to_led_control_port_slave_write),         //                                           .write
		.dma_ssram_to_led_control_port_slave_readdata      (mm_interconnect_0_dma_ssram_to_led_control_port_slave_readdata),      //                                           .readdata
		.dma_ssram_to_led_control_port_slave_writedata     (mm_interconnect_0_dma_ssram_to_led_control_port_slave_writedata),     //                                           .writedata
		.dma_ssram_to_led_control_port_slave_chipselect    (mm_interconnect_0_dma_ssram_to_led_control_port_slave_chipselect),    //                                           .chipselect
		.led_fifo_in_address                               (mm_interconnect_0_led_fifo_in_address),                               //                                led_fifo_in.address
		.led_fifo_in_write                                 (mm_interconnect_0_led_fifo_in_write),                                 //                                           .write
		.led_fifo_in_writedata                             (mm_interconnect_0_led_fifo_in_writedata),                             //                                           .writedata
		.led_fifo_in_waitrequest                           (mm_interconnect_0_led_fifo_in_waitrequest),                           //                                           .waitrequest
		.led_out_led_address                               (mm_interconnect_0_led_out_led_address),                               //                                led_out_led.address
		.led_out_led_write                                 (mm_interconnect_0_led_out_led_write),                                 //                                           .write
		.led_out_led_read                                  (mm_interconnect_0_led_out_led_read),                                  //                                           .read
		.led_out_led_readdata                              (mm_interconnect_0_led_out_led_readdata),                              //                                           .readdata
		.led_out_led_writedata                             (mm_interconnect_0_led_out_led_writedata),                             //                                           .writedata
		.test_mem_s1_address                               (mm_interconnect_0_test_mem_s1_address),                               //                                test_mem_s1.address
		.test_mem_s1_write                                 (mm_interconnect_0_test_mem_s1_write),                                 //                                           .write
		.test_mem_s1_readdata                              (mm_interconnect_0_test_mem_s1_readdata),                              //                                           .readdata
		.test_mem_s1_writedata                             (mm_interconnect_0_test_mem_s1_writedata),                             //                                           .writedata
		.test_mem_s1_byteenable                            (mm_interconnect_0_test_mem_s1_byteenable),                            //                                           .byteenable
		.test_mem_s1_chipselect                            (mm_interconnect_0_test_mem_s1_chipselect),                            //                                           .chipselect
		.test_mem_s1_clken                                 (mm_interconnect_0_test_mem_s1_clken)                                  //                                           .clken
	);

	sm_transfer_system_mm_interconnect_1 mm_interconnect_1 (
		.pll_outclk0_clk                                       (pll_outclk0_clk),                               //                                     pll_outclk0.clk
		.dma_source_to_ssram_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                // dma_source_to_ssram_reset_reset_bridge_in_reset.reset
		.dma_source_to_ssram_read_master_address               (dma_source_to_ssram_read_master_address),       //                 dma_source_to_ssram_read_master.address
		.dma_source_to_ssram_read_master_waitrequest           (dma_source_to_ssram_read_master_waitrequest),   //                                                .waitrequest
		.dma_source_to_ssram_read_master_chipselect            (dma_source_to_ssram_read_master_chipselect),    //                                                .chipselect
		.dma_source_to_ssram_read_master_read                  (~dma_source_to_ssram_read_master_read),         //                                                .read
		.dma_source_to_ssram_read_master_readdata              (dma_source_to_ssram_read_master_readdata),      //                                                .readdata
		.dma_source_to_ssram_read_master_readdatavalid         (dma_source_to_ssram_read_master_readdatavalid), //                                                .readdatavalid
		.source_s1_address                                     (mm_interconnect_1_source_s1_address),           //                                       source_s1.address
		.source_s1_write                                       (mm_interconnect_1_source_s1_write),             //                                                .write
		.source_s1_readdata                                    (mm_interconnect_1_source_s1_readdata),          //                                                .readdata
		.source_s1_writedata                                   (mm_interconnect_1_source_s1_writedata),         //                                                .writedata
		.source_s1_byteenable                                  (mm_interconnect_1_source_s1_byteenable),        //                                                .byteenable
		.source_s1_chipselect                                  (mm_interconnect_1_source_s1_chipselect),        //                                                .chipselect
		.source_s1_clken                                       (mm_interconnect_1_source_s1_clken),             //                                                .clken
		.source_s1_debugaccess                                 (mm_interconnect_1_source_s1_debugaccess)        //                                                .debugaccess
	);

	sm_transfer_system_mm_interconnect_2 mm_interconnect_2 (
		.pll_outclk0_clk                                    (pll_outclk0_clk),                                     //                                  pll_outclk0.clk
		.dma_ssram_to_led_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                      // dma_ssram_to_led_reset_reset_bridge_in_reset.reset
		.dma_source_to_ssram_write_master_address           (dma_source_to_ssram_write_master_address),            //             dma_source_to_ssram_write_master.address
		.dma_source_to_ssram_write_master_waitrequest       (dma_source_to_ssram_write_master_waitrequest),        //                                             .waitrequest
		.dma_source_to_ssram_write_master_byteenable        (dma_source_to_ssram_write_master_byteenable),         //                                             .byteenable
		.dma_source_to_ssram_write_master_chipselect        (dma_source_to_ssram_write_master_chipselect),         //                                             .chipselect
		.dma_source_to_ssram_write_master_write             (~dma_source_to_ssram_write_master_write),             //                                             .write
		.dma_source_to_ssram_write_master_writedata         (dma_source_to_ssram_write_master_writedata),          //                                             .writedata
		.dma_ssram_to_led_read_master_address               (dma_ssram_to_led_read_master_address),                //                 dma_ssram_to_led_read_master.address
		.dma_ssram_to_led_read_master_waitrequest           (dma_ssram_to_led_read_master_waitrequest),            //                                             .waitrequest
		.dma_ssram_to_led_read_master_chipselect            (dma_ssram_to_led_read_master_chipselect),             //                                             .chipselect
		.dma_ssram_to_led_read_master_read                  (~dma_ssram_to_led_read_master_read),                  //                                             .read
		.dma_ssram_to_led_read_master_readdata              (dma_ssram_to_led_read_master_readdata),               //                                             .readdata
		.dma_ssram_to_led_read_master_readdatavalid         (dma_ssram_to_led_read_master_readdatavalid),          //                                             .readdatavalid
		.sram_controller_uas_address                        (mm_interconnect_2_sram_controller_uas_address),       //                          sram_controller_uas.address
		.sram_controller_uas_write                          (mm_interconnect_2_sram_controller_uas_write),         //                                             .write
		.sram_controller_uas_read                           (mm_interconnect_2_sram_controller_uas_read),          //                                             .read
		.sram_controller_uas_readdata                       (mm_interconnect_2_sram_controller_uas_readdata),      //                                             .readdata
		.sram_controller_uas_writedata                      (mm_interconnect_2_sram_controller_uas_writedata),     //                                             .writedata
		.sram_controller_uas_burstcount                     (mm_interconnect_2_sram_controller_uas_burstcount),    //                                             .burstcount
		.sram_controller_uas_byteenable                     (mm_interconnect_2_sram_controller_uas_byteenable),    //                                             .byteenable
		.sram_controller_uas_readdatavalid                  (mm_interconnect_2_sram_controller_uas_readdatavalid), //                                             .readdatavalid
		.sram_controller_uas_waitrequest                    (mm_interconnect_2_sram_controller_uas_waitrequest),   //                                             .waitrequest
		.sram_controller_uas_lock                           (mm_interconnect_2_sram_controller_uas_lock),          //                                             .lock
		.sram_controller_uas_debugaccess                    (mm_interconnect_2_sram_controller_uas_debugaccess)    //                                             .debugaccess
	);

	sm_transfer_system_avalon_st_adapter #(
		.inBitsPerSymbol (32),
		.inUsePackets    (0),
		.inDataWidth     (32),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (32),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk   (pll_outclk0_clk),                // in_clk_0.clk
		.in_rst_0_reset (rst_controller_reset_out_reset), // in_rst_0.reset
		.in_0_data      (led_fifo_out_data),              //     in_0.data
		.in_0_valid     (led_fifo_out_valid),             //         .valid
		.in_0_ready     (led_fifo_out_ready),             //         .ready
		.out_0_data     (avalon_st_adapter_out_0_data),   //    out_0.data
		.out_0_valid    (avalon_st_adapter_out_0_valid),  //         .valid
		.out_0_ready    (avalon_st_adapter_out_0_ready)   //         .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_debounce_button_qual_reset), // reset_in0.reset
		.reset_in1      (j2a_master_master_reset_reset),    // reset_in1.reset
		.clk            (pll_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                 // (terminated)
		.reset_req_in0  (1'b0),                             // (terminated)
		.reset_req_in1  (1'b0),                             // (terminated)
		.reset_in2      (1'b0),                             // (terminated)
		.reset_req_in2  (1'b0),                             // (terminated)
		.reset_in3      (1'b0),                             // (terminated)
		.reset_req_in3  (1'b0),                             // (terminated)
		.reset_in4      (1'b0),                             // (terminated)
		.reset_req_in4  (1'b0),                             // (terminated)
		.reset_in5      (1'b0),                             // (terminated)
		.reset_req_in5  (1'b0),                             // (terminated)
		.reset_in6      (1'b0),                             // (terminated)
		.reset_req_in6  (1'b0),                             // (terminated)
		.reset_in7      (1'b0),                             // (terminated)
		.reset_req_in7  (1'b0),                             // (terminated)
		.reset_in8      (1'b0),                             // (terminated)
		.reset_req_in8  (1'b0),                             // (terminated)
		.reset_in9      (1'b0),                             // (terminated)
		.reset_req_in9  (1'b0),                             // (terminated)
		.reset_in10     (1'b0),                             // (terminated)
		.reset_req_in10 (1'b0),                             // (terminated)
		.reset_in11     (1'b0),                             // (terminated)
		.reset_req_in11 (1'b0),                             // (terminated)
		.reset_in12     (1'b0),                             // (terminated)
		.reset_req_in12 (1'b0),                             // (terminated)
		.reset_in13     (1'b0),                             // (terminated)
		.reset_req_in13 (1'b0),                             // (terminated)
		.reset_in14     (1'b0),                             // (terminated)
		.reset_req_in14 (1'b0),                             // (terminated)
		.reset_in15     (1'b0),                             // (terminated)
		.reset_req_in15 (1'b0)                              // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (j2a_master_master_reset_reset),      // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
