
module unnamed (
	clk_clk,
	pio_0_external_connection_export,
	pio_1_external_connection_export);	

	input		clk_clk;
	input		pio_0_external_connection_export;
	output		pio_1_external_connection_export;
endmodule
