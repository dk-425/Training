
module unsaved (
	blink_0_avalon_slave_0_beginbursttransfer,
	blink_0_avalon_slave_0_writeresponsevalid_n);	

	input		blink_0_avalon_slave_0_beginbursttransfer;
	output		blink_0_avalon_slave_0_writeresponsevalid_n;
endmodule
