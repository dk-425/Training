`timescale 1ns / 1ps

module axistb(

    );
    reg clk;
    reg reset_n;
    reg [7:0] s_tdata;
    reg s_tlast;
    reg s_tvalid;  
    reg m_tready;
    wire s_tready;   
    wire [7:0] m_tdata;
    wire m_tvalid;
      
    // Instantiating
   axis_reg #(
        .N(8)
    ) dut (
        .clk(clk),
        .reset_n(reset_n),
        .s_tdata(s_tdata),
        .s_tvalid(s_tvalid),
        .s_tready(s_tready),
        .s_tlast(s_tlast),
        .m_tdata(m_tdata),
        .m_tvalid(m_tvalid),
        .m_tready(m_tready)
    );
   /*  design_1_wrapper uut
   (.clk_0(clk),
    .m_0_tdata(m_tdata),
    .m_0_tvalid(m_tvalid),
    .reset_n_0(reset_n),
    .s_0_tdata(s_tdata),
    .s_0_tlast(s_tlast),
    .s_0_tready(s_tready),
    .s_0_tvalid(s_tvalid),
    .m_0_tready(m_tready));
    */
    // Clock generation
    always #5 clk = ~clk;
    
    initial begin
        // Initialize inputs
        clk = 0;
        reset_n = 1;
        s_tdata = 8'h00;
        s_tvalid = 0;
        
        
        // Apply reset
        reset_n <= 0;
        #10;
        reset_n <= 1;
        m_tready<=1;
        
        
        // Send data and wait for it to be accepted
        s_tdata <= 8'b01101000;
        s_tlast <= 1'b1;
        
        #1
        
        s_tvalid <= 1;
        #10;
        s_tvalid <= 0;
        #40
        m_tready<=0;
        #5
        // Finish simulation
        $finish;
    end

endmodule
